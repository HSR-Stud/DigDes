resize(a, y'length) --auf Laenge von y
resize(b, 8) -- auf 8bit
