component <COMPONENT_NAME>
	port(
		{<PORT_NAME>: <mode> <type>;});
end component;
