signal <sig_name> {, <sig_name>}: <type>;
